
module Fifo #(parameter DATA_WIDTH = 8,
              parameter DEPTH = 16)
             (input clk,                          // clock, active when posedge
              input reset,                        // synchronous reset; active high
              input rd_enable,
              input wr_enable,                    // if the data_in is passenger, enable = 1; if the data_in is luggage, enable = 0
              input [DATA_WIDTH-1:0] data_in,
              output reg [DATA_WIDTH-1:0] data_out,
              output reg full, empty);
    localparam PTR_WIDTH = $clog2(DEPTH);

    reg [DATA_WIDTH-1:0] fifo[DEPTH-1:0];
    reg [PTR_WIDTH-1:0] write_ptr = 0, read_ptr = 0; // pointers to the stack


    always@(posedge clk) begin
        if (reset) begin
            write_ptr <= 0;
            read_ptr  <= 0;
        end
        else begin
            if (!full && wr_enable) begin
                fifo[write_ptr] <= data_in;
                write_ptr       <= ((write_ptr + 1) % DEPTH);
            end
            if (!empty && rd_enable) begin
                data_out <= fifo[read_ptr];
                read_ptr <= ((read_ptr + 1) % DEPTH);
            end
        end
    end
    assign full  = (((write_ptr + 1) % DEPTH) == read_ptr);
    assign empty = (write_ptr == read_ptr);
endmodule


// // testbench
// module Fifo_tb;
//     reg clk, rst, wr_en, rd_en;
//     reg [7:0] data_in;
//     wire [7:0] data_out;
//     wire full, empty;

//     Fifo #(8, 16) fifo(.clk(clk), .reset(rst),
//     .wr_enable(en),
//     .rd_enable(en),
//     .data_in(data_in),
//     .data_out(data_out),
//     .full(full),
//     .empty(empty));

//     initial begin
//         clk = 0;
//         forever #5 clk = ~clk;  // Clock generation
//     end

//     initial begin
//         rst = 1;
//         wr_en = 0;
//         rd_en = 0;
//         data_in = 8'h0;
//         #10 rst = 0;  // Release reset

//         // Begin test sequence
//         wr_en = 1;
//         data_in = 8'hA; #10;
//         data_in = 8'hB; #10;
//         data_in = 8'hC; #10;
//         data_in = 8'hD; #10;


//         // Testing ENABLE = 0
//         wr_en = 0;
//         rd_en = 1;
//         data_in = 8'h1; #10;
//         data_in = 8'h2; #10;
//         data_in = 8'h3; #10;


//         #10 $display("time = %d, clk = %d, data_out = %h", $time, clk, data_out);
//         #10 $display("time = %d, clk = %d, data_out = %h", $time, clk, data_out);
//         #10 $display("time = %d, clk = %d, data_out = %h", $time, clk, data_out);
//         #10 $display("time = %d, clk = %d, data_out = %h", $time, clk, data_out);
//         #10 $display("time = %d, clk = %d, data_out = %h", $time, clk, data_out);

//         $finish;  // End simulation
//     end
// endmodule
